module dec16to40(input [15:0] select,output reg [39:0] decout);
	always@(select)
	begin
	case(select)
	16'b0000000000000000:decout=40'b0000000000000000000000000000000000000001;
	16'b0000000000000001:decout=40'b0000000000000000000000000000000000000010;
	16'b0000000000000010:decout=40'b0000000000000000000000000000000000000100;
	16'b0000000000000011:decout=40'b0000000000000000000000000000000000001000;
	16'b0000000000000100:decout=40'b0000000000000000000000000000000000010000;
	16'b0000000000000101:decout=40'b0000000000000000000000000000000000100000;
	16'b0000000000000110:decout=40'b0000000000000000000000000000000001000000;
	16'b0000000000000111:decout=40'b0000000000000000000000000000000010000000;
	16'b0000000000001000:decout=40'b0000000000000000000000000000000100000000;
	16'b0000000000001001:decout=40'b0000000000000000000000000000001000000000;
	16'b0000000000001010:decout=40'b0000000000000000000000000000010000000000;
	16'b0000000000001011:decout=40'b0000000000000000000000000000100000000000;
	16'b0000000000001100:decout=40'b0000000000000000000000000001000000000000;
	16'b0000000000001101:decout=40'b0000000000000000000000000010000000000000;
	16'b0000000000001110:decout=40'b0000000000000000000000000100000000000000;
	16'b0000000000001111:decout=40'b0000000000000000000000001000000000000000;
	16'b0000000000010000:decout=40'b0000000000000000000000010000000000000000;
	16'b0000000000010001:decout=40'b0000000000000000000000100000000000000000;
	16'b0000000000010010:decout=40'b0000000000000000000001000000000000000000;
	16'b0000000000010011:decout=40'b0000000000000000000010000000000000000000;
	16'b0000000000010100:decout=40'b0000000000000000000100000000000000000000;
	16'b0000000000010101:decout=40'b0000000000000000001000000000000000000000;
	16'b0000000000010110:decout=40'b0000000000000000010000000000000000000000;
	16'b0000000000010111:decout=40'b0000000000000000100000000000000000000000;
	16'b0000000000011000:decout=40'b0000000000000001000000000000000000000000;
	16'b0000000000011001:decout=40'b0000000000000010000000000000000000000000;
	16'b0000000000011010:decout=40'b0000000000000100000000000000000000000000;
	16'b0000000000011011:decout=40'b0000000000001000000000000000000000000000;
	16'b0000000000011100:decout=40'b0000000000010000000000000000000000000000;
	16'b0000000000011101:decout=40'b0000000000100000000000000000000000000000;
	16'b0000000000011110:decout=40'b0000000001000000000000000000000000000000;
	16'b0000000000011111:decout=40'b0000000010000000000000000000000000000000;
	16'b0000000000100000:decout=40'b0000000100000000000000000000000000000000;
	16'b0000000000100001:decout=40'b0000001000000000000000000000000000000000;
	16'b0000000000100010:decout=40'b0000010000000000000000000000000000000000;
	16'b0000000000100011:decout=40'b0000100000000000000000000000000000000000;
	16'b0000000000100100:decout=40'b0001000000000000000000000000000000000000;
	16'b0000000000100101:decout=40'b0010000000000000000000000000000000000000;
	16'b0000000000100110:decout=40'b0100000000000000000000000000000000000000;
	16'b0000000000100111:decout=40'b1000000000000000000000000000000000000000;
	endcase
	end
endmodule